/filespace/k/krasselt/ECE755/ECE755_SP25_Project/Milestone_4/asap7sc7p5t_28/techlef_misc/asap7_tech_4x_201209.lef