/filespace/k/krasselt/ECE755/ECE755_SP25_Project/Milestone_4/asap7sc7p5t_28/LEF/scaled/asap7sc7p5t_28_R_4x_220121a.lef